`timescale 1ns / 1ps
// =============================================================================
//  Program : distri_ram.v
//  Author  : Dong-Fong Syu
//  Date    : Feb/01/2018
// -----------------------------------------------------------------------------
//  Description:
//  This is the Distributed RAM module for the Aquila core (A RISC-V core).
// -----------------------------------------------------------------------------
//  Revision information:
//
//  None.
// -----------------------------------------------------------------------------
//  License information:
//
//  This software is released under the BSD-3-Clause Licence,
//  see https://opensource.org/licenses/BSD-3-Clause for details.
//  In the following license statements, "software" refers to the
//  "source code" of the complete hardware/software system.
//
//  Copyright 2019,
//                    Embedded Intelligent Systems Lab (EISL)
//                    Deparment of Computer Science
//                    National Chiao Tung Uniersity
//                    Hsinchu, Taiwan.s
//
//  All rights reserved.
//
//  Redistribution and use in source and binary forms, with or without
//  modification, are permitted provided that the following conditions are met:
//
//  1. Redistributions of source code must retain the above copyright notice,
//     this list of conditions and the following disclaimer.
//
//  2. Redistributions in binary form must reproduce the above copyright notice,
//     this list of conditions and the following disclaimer in the documentation
//     and/or other materials provided with the distribution.
//
//  3. Neither the name of the copyright holder nor the names of its contributors
//     may be used to endorse or promote products derived from this software
//     without specific prior written permission.
//
//  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
//  AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
//  IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
//  ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
//  LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
//  CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
//  SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
//  INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
//  CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
//  ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
//  POSSIBILITY OF SUCH DAMAGE.
// =============================================================================

module distri_ram_dp
#(parameter ENTRY_NUM = 32,
  parameter XLEN = 32,
  parameter AWDTH = $clog2(ENTRY_NUM))
(
    input                clk_i,
    input  [XLEN-1 : 0]  data_i,
    input                we_i,
    input  [AWDTH-1 : 0] write_addr_i,

    input  [AWDTH-1 : 0] a_read_addr_i,
    output [XLEN-1 : 0]  a_data_o,

    input  [AWDTH-1 : 0] b_read_addr_i,
    output [XLEN-1 : 0]  b_data_o
);

reg [XLEN-1 : 0] RAM[ENTRY_NUM-1 : 0];
integer i;

assign a_data_o = RAM[a_read_addr_i];
assign b_data_o = RAM[b_read_addr_i];

initial
begin
    for (i = 0; i < ENTRY_NUM; i = i + 1)
        RAM[i] <= 0;
end

always @(posedge clk_i)
begin
    if (we_i)
    begin
        RAM[write_addr_i] <= data_i;
    end
end



endmodule
