`timescale 1ns / 1ps
// =============================================================================
//  Program : bram_dp_L2.v
//  Author  : Lin-en Yen
//  Date    : Apr/1/2024
// -----------------------------------------------------------------------------
//  Description:
//  This module synthesizes an SRAM with output 'data_o' in latch mode.
//  when 'we_i' is enabled, 'data_i' will be feed to 'data_o' before the
//  next clock rising edge.
// -----------------------------------------------------------------------------
//  Revision information:
//
//  None.
// -----------------------------------------------------------------------------
//  License information:
//
//  This software is released under the BSD-3-Clause Licence,
//  see https://opensource.org/licenses/BSD-3-Clause for details.
//  In the following license statements, "software" refers to the
//  "source code" of the complete hardware/software system.
//
//  Copyright 2023,
//                    Embedded Intelligent Systems Lab (EISL)
//                    Deparment of Computer Science
//                    National Yang Ming Chiao Tung Uniersity (NYCU)
//                    Hsinchu, Taiwan.
//
//  All rights reserved.
//
//  Redistribution and use in source and binary forms, with or without
//  modification, are permitted provided that the following conditions are met:
//
//  1. Redistributions of source code must retain the above copyright notice,
//     this list of conditions and the following disclaimer.
//
//  2. Redistributions in binary form must reproduce the above copyright notice,
//     this list of conditions and the following disclaimer in the documentation
//     and/or other materials provided with the distribution.
//
//  3. Neither the name of the copyright holder nor the names of its contributors
//     may be used to endorse or promote products derived from this software
//     without specific prior written permission.
//
//  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
//  AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
//  IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
//  ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
//  LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
//  CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
//  SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
//  INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
//  CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
//  ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
//  POSSIBILITY OF SUCH DAMAGE.
// =============================================================================

module bram_dp
#(parameter DATA_WIDTH = 32, N_ENTRIES = 128)
(
    input                           clk_i,
    input                           en_i,
    input                           a_we_i,
    input  [$clog2(N_ENTRIES)-1: 0] a_addr_i,
    input  [DATA_WIDTH-1: 0]        a_data_i,
    output reg [DATA_WIDTH-1: 0]    a_data_o,

    input                           b_we_i,
    input  [$clog2(N_ENTRIES)-1: 0] b_addr_i,
    input  [DATA_WIDTH-1: 0]        b_data_i,
    output reg [DATA_WIDTH-1: 0]    b_data_o
);

reg [DATA_WIDTH-1 : 0] RAM [N_ENTRIES-1: 0];

always @(posedge clk_i)
begin
    if (en_i)
    begin
        if (a_we_i)
        begin
            RAM[a_addr_i] <= a_data_i;
            a_data_o <= a_data_i;
        end
        else
            a_data_o <= RAM[a_addr_i];
    end
end

always @(posedge clk_i)
begin
    if (en_i)
    begin
        if (b_we_i)
        begin
            RAM[b_addr_i] <= b_data_i;
            b_data_o <= b_data_i;
        end
        else
            b_data_o <= RAM[b_addr_i];
    end
end

endmodule
